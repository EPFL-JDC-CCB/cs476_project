`default_nettype none 
module charRom ( input wire        clock,
                 input wire [9:0] address,
                 output reg [7:0]  data);

  always @(posedge clock)
  begin
    case (address)
      10'h008 : data <= 8'h7E;
      10'h009 : data <= 8'h81;
      10'h00A : data <= 8'hA5;
      10'h00B : data <= 8'h81;
      10'h00C : data <= 8'hBD;
      10'h00D : data <= 8'h99;
      10'h00E : data <= 8'h81;
      10'h00F : data <= 8'h7E;
      10'h010 : data <= 8'h7E;
      10'h011 : data <= 8'hFF;
      10'h012 : data <= 8'hDB;
      10'h013 : data <= 8'hFF;
      10'h014 : data <= 8'hC3;
      10'h015 : data <= 8'hE7;
      10'h016 : data <= 8'hFF;
      10'h017 : data <= 8'h7E;
      10'h018 : data <= 8'h44;
      10'h019 : data <= 8'hEE;
      10'h01A : data <= 8'hFE;
      10'h01B : data <= 8'hFE;
      10'h01C : data <= 8'h7C;
      10'h01D : data <= 8'h38;
      10'h01E : data <= 8'h10;
      10'h020 : data <= 8'h10;
      10'h021 : data <= 8'h38;
      10'h022 : data <= 8'h7C;
      10'h023 : data <= 8'hFE;
      10'h024 : data <= 8'h7C;
      10'h025 : data <= 8'h38;
      10'h026 : data <= 8'h10;
      10'h028 : data <= 8'h18;
      10'h029 : data <= 8'h3C;
      10'h02A : data <= 8'hDB;
      10'h02B : data <= 8'hFF;
      10'h02C : data <= 8'hDB;
      10'h02D : data <= 8'h18;
      10'h02E : data <= 8'h3C;
      10'h030 : data <= 8'h18;
      10'h031 : data <= 8'h3C;
      10'h032 : data <= 8'h7E;
      10'h033 : data <= 8'hFF;
      10'h034 : data <= 8'h7E;
      10'h035 : data <= 8'h18;
      10'h036 : data <= 8'h3C;
      10'h03A : data <= 8'h3C;
      10'h03B : data <= 8'h3C;
      10'h03C : data <= 8'h3C;
      10'h03D : data <= 8'h3C;
      10'h040 : data <= 8'hFF;
      10'h041 : data <= 8'hFF;
      10'h042 : data <= 8'hC3;
      10'h043 : data <= 8'hC3;
      10'h044 : data <= 8'hC3;
      10'h045 : data <= 8'hC3;
      10'h046 : data <= 8'hFF;
      10'h047 : data <= 8'hFF;
      10'h049 : data <= 8'h7E;
      10'h04A : data <= 8'h42;
      10'h04B : data <= 8'h42;
      10'h04C : data <= 8'h42;
      10'h04D : data <= 8'h42;
      10'h04E : data <= 8'h7E;
      10'h050 : data <= 8'hFF;
      10'h051 : data <= 8'h81;
      10'h052 : data <= 8'hBD;
      10'h053 : data <= 8'hBD;
      10'h054 : data <= 8'hBD;
      10'h055 : data <= 8'hBD;
      10'h056 : data <= 8'h81;
      10'h057 : data <= 8'hFF;
      10'h058 : data <= 8'h0F;
      10'h059 : data <= 8'h07;
      10'h05A : data <= 8'h07;
      10'h05B : data <= 8'h7D;
      10'h05C : data <= 8'hCC;
      10'h05D : data <= 8'hCC;
      10'h05E : data <= 8'hCC;
      10'h05F : data <= 8'h78;
      10'h060 : data <= 8'h78;
      10'h061 : data <= 8'hCC;
      10'h062 : data <= 8'hCC;
      10'h063 : data <= 8'hCC;
      10'h064 : data <= 8'h78;
      10'h065 : data <= 8'h30;
      10'h066 : data <= 8'hFC;
      10'h067 : data <= 8'h30;
      10'h068 : data <= 8'h1F;
      10'h069 : data <= 8'h33;
      10'h06A : data <= 8'h3F;
      10'h06B : data <= 8'h30;
      10'h06C : data <= 8'h30;
      10'h06D : data <= 8'h70;
      10'h06E : data <= 8'hF0;
      10'h06F : data <= 8'hE0;
      10'h070 : data <= 8'h3F;
      10'h071 : data <= 8'h63;
      10'h072 : data <= 8'h7F;
      10'h073 : data <= 8'h63;
      10'h074 : data <= 8'h63;
      10'h075 : data <= 8'h67;
      10'h076 : data <= 8'hE6;
      10'h077 : data <= 8'hC0;
      10'h078 : data <= 8'hDB;
      10'h079 : data <= 8'hDB;
      10'h07A : data <= 8'h3C;
      10'h07B : data <= 8'hE7;
      10'h07C : data <= 8'hE7;
      10'h07D : data <= 8'h3C;
      10'h07E : data <= 8'hDB;
      10'h07F : data <= 8'hDB;
      10'h080 : data <= 8'hC0;
      10'h081 : data <= 8'hF0;
      10'h082 : data <= 8'hF8;
      10'h083 : data <= 8'hFE;
      10'h084 : data <= 8'hF8;
      10'h085 : data <= 8'hF0;
      10'h086 : data <= 8'hC0;
      10'h088 : data <= 8'h06;
      10'h089 : data <= 8'h1E;
      10'h08A : data <= 8'h3E;
      10'h08B : data <= 8'hFE;
      10'h08C : data <= 8'h3E;
      10'h08D : data <= 8'h1E;
      10'h08E : data <= 8'h06;
      10'h090 : data <= 8'h30;
      10'h091 : data <= 8'h78;
      10'h092 : data <= 8'hFC;
      10'h093 : data <= 8'h30;
      10'h094 : data <= 8'h30;
      10'h095 : data <= 8'hFC;
      10'h096 : data <= 8'h78;
      10'h097 : data <= 8'h30;
      10'h098 : data <= 8'h6C;
      10'h099 : data <= 8'h6C;
      10'h09A : data <= 8'h6C;
      10'h09B : data <= 8'h6C;
      10'h09C : data <= 8'h6C;
      10'h09E : data <= 8'h6C;
      10'h0A0 : data <= 8'h7F;
      10'h0A1 : data <= 8'hDB;
      10'h0A2 : data <= 8'hDB;
      10'h0A3 : data <= 8'hDB;
      10'h0A4 : data <= 8'h7B;
      10'h0A5 : data <= 8'h1B;
      10'h0A6 : data <= 8'h1B;
      10'h0A8 : data <= 8'h3C;
      10'h0A9 : data <= 8'h60;
      10'h0AA : data <= 8'h3C;
      10'h0AB : data <= 8'h66;
      10'h0AC : data <= 8'h66;
      10'h0AD : data <= 8'h3C;
      10'h0AE : data <= 8'h06;
      10'h0AF : data <= 8'h3C;
      10'h0B4 : data <= 8'hFE;
      10'h0B5 : data <= 8'hFE;
      10'h0B6 : data <= 8'hFE;
      10'h0B8 : data <= 8'h18;
      10'h0B9 : data <= 8'h3C;
      10'h0BA : data <= 8'h7E;
      10'h0BB : data <= 8'h18;
      10'h0BC : data <= 8'h7E;
      10'h0BD : data <= 8'h3C;
      10'h0BE : data <= 8'h18;
      10'h0BF : data <= 8'h7E;
      10'h0C0 : data <= 8'h30;
      10'h0C1 : data <= 8'h78;
      10'h0C2 : data <= 8'hFC;
      10'h0C3 : data <= 8'h30;
      10'h0C4 : data <= 8'h30;
      10'h0C5 : data <= 8'h30;
      10'h0C6 : data <= 8'h30;
      10'h0C8 : data <= 8'h30;
      10'h0C9 : data <= 8'h30;
      10'h0CA : data <= 8'h30;
      10'h0CB : data <= 8'h30;
      10'h0CC : data <= 8'hFC;
      10'h0CD : data <= 8'h78;
      10'h0CE : data <= 8'h30;
      10'h0D1 : data <= 8'h08;
      10'h0D2 : data <= 8'h0C;
      10'h0D3 : data <= 8'hFE;
      10'h0D4 : data <= 8'h0C;
      10'h0D5 : data <= 8'h08;
      10'h0D9 : data <= 8'h20;
      10'h0DA : data <= 8'h60;
      10'h0DB : data <= 8'hFE;
      10'h0DC : data <= 8'h60;
      10'h0DD : data <= 8'h20;
      10'h0E2 : data <= 8'hC0;
      10'h0E3 : data <= 8'hC0;
      10'h0E4 : data <= 8'hFE;
      10'h0E9 : data <= 8'h24;
      10'h0EA : data <= 8'h42;
      10'h0EB : data <= 8'hFF;
      10'h0EC : data <= 8'h42;
      10'h0ED : data <= 8'h24;
      10'h0F1 : data <= 8'h10;
      10'h0F2 : data <= 8'h38;
      10'h0F3 : data <= 8'h7C;
      10'h0F4 : data <= 8'hFE;
      10'h0F5 : data <= 8'hFE;
      10'h0F9 : data <= 8'hFE;
      10'h0FA : data <= 8'hFE;
      10'h0FB : data <= 8'h7C;
      10'h0FC : data <= 8'h38;
      10'h0FD : data <= 8'h10;
      10'h108 : data <= 8'h18;
      10'h109 : data <= 8'h18;
      10'h10A : data <= 8'h18;
      10'h10B : data <= 8'h18;
      10'h10C : data <= 8'h18;
      10'h10E : data <= 8'h18;
      10'h110 : data <= 8'hCC;
      10'h111 : data <= 8'hCC;
      10'h112 : data <= 8'hCC;
      10'h118 : data <= 8'h36;
      10'h119 : data <= 8'h6C;
      10'h11A : data <= 8'hFE;
      10'h11B : data <= 8'h6C;
      10'h11C : data <= 8'hFE;
      10'h11D : data <= 8'h6C;
      10'h11E : data <= 8'hD8;
      10'h120 : data <= 8'h18;
      10'h121 : data <= 8'h7E;
      10'h122 : data <= 8'hC0;
      10'h123 : data <= 8'h7C;
      10'h124 : data <= 8'h06;
      10'h125 : data <= 8'hFC;
      10'h126 : data <= 8'h30;
      10'h128 : data <= 8'hC2;
      10'h129 : data <= 8'hC6;
      10'h12A : data <= 8'h0C;
      10'h12B : data <= 8'h18;
      10'h12C : data <= 8'h30;
      10'h12D : data <= 8'h66;
      10'h12E : data <= 8'hC6;
      10'h130 : data <= 8'h38;
      10'h131 : data <= 8'h6C;
      10'h132 : data <= 8'h38;
      10'h133 : data <= 8'h70;
      10'h134 : data <= 8'hDE;
      10'h135 : data <= 8'hCC;
      10'h136 : data <= 8'h76;
      10'h138 : data <= 8'h30;
      10'h139 : data <= 8'h30;
      10'h13A : data <= 8'h60;
      10'h140 : data <= 8'h0C;
      10'h141 : data <= 8'h18;
      10'h142 : data <= 8'h30;
      10'h143 : data <= 8'h30;
      10'h144 : data <= 8'h30;
      10'h145 : data <= 8'h18;
      10'h146 : data <= 8'h0C;
      10'h148 : data <= 8'h30;
      10'h149 : data <= 8'h18;
      10'h14A : data <= 8'h0C;
      10'h14B : data <= 8'h0C;
      10'h14C : data <= 8'h0C;
      10'h14D : data <= 8'h18;
      10'h14E : data <= 8'h30;
      10'h151 : data <= 8'h6C;
      10'h152 : data <= 8'h38;
      10'h153 : data <= 8'hFE;
      10'h154 : data <= 8'h38;
      10'h155 : data <= 8'h6C;
      10'h159 : data <= 8'h18;
      10'h15A : data <= 8'h18;
      10'h15B : data <= 8'h7E;
      10'h15C : data <= 8'h18;
      10'h15D : data <= 8'h18;
      10'h165 : data <= 8'h18;
      10'h166 : data <= 8'h18;
      10'h167 : data <= 8'h30;
      10'h16B : data <= 8'h7E;
      10'h175 : data <= 8'h18;
      10'h176 : data <= 8'h18;
      10'h178 : data <= 8'h02;
      10'h179 : data <= 8'h06;
      10'h17A : data <= 8'h0C;
      10'h17B : data <= 8'h18;
      10'h17C : data <= 8'h30;
      10'h17D : data <= 8'h60;
      10'h17E : data <= 8'hC0;
      10'h180 : data <= 8'h7C;
      10'h181 : data <= 8'hCE;
      10'h182 : data <= 8'hDE;
      10'h183 : data <= 8'hF6;
      10'h184 : data <= 8'hE6;
      10'h185 : data <= 8'hC6;
      10'h186 : data <= 8'h7C;
      10'h188 : data <= 8'h18;
      10'h189 : data <= 8'h38;
      10'h18A : data <= 8'h18;
      10'h18B : data <= 8'h18;
      10'h18C : data <= 8'h18;
      10'h18D : data <= 8'h18;
      10'h18E : data <= 8'h7E;
      10'h190 : data <= 8'h7C;
      10'h191 : data <= 8'hC6;
      10'h192 : data <= 8'h06;
      10'h193 : data <= 8'h1C;
      10'h194 : data <= 8'h70;
      10'h195 : data <= 8'hC6;
      10'h196 : data <= 8'hFE;
      10'h198 : data <= 8'h7C;
      10'h199 : data <= 8'hC6;
      10'h19A : data <= 8'h06;
      10'h19B : data <= 8'h1C;
      10'h19C : data <= 8'h06;
      10'h19D : data <= 8'hC6;
      10'h19E : data <= 8'h7C;
      10'h1A0 : data <= 8'h1C;
      10'h1A1 : data <= 8'h3C;
      10'h1A2 : data <= 8'h6C;
      10'h1A3 : data <= 8'hCC;
      10'h1A4 : data <= 8'hFE;
      10'h1A5 : data <= 8'h0C;
      10'h1A6 : data <= 8'h0C;
      10'h1A8 : data <= 8'hFE;
      10'h1A9 : data <= 8'hC0;
      10'h1AA : data <= 8'hFC;
      10'h1AB : data <= 8'h06;
      10'h1AC : data <= 8'h06;
      10'h1AD : data <= 8'hC6;
      10'h1AE : data <= 8'h7C;
      10'h1B0 : data <= 8'h3C;
      10'h1B1 : data <= 8'h60;
      10'h1B2 : data <= 8'hC0;
      10'h1B3 : data <= 8'hFC;
      10'h1B4 : data <= 8'hC6;
      10'h1B5 : data <= 8'hC6;
      10'h1B6 : data <= 8'h7C;
      10'h1B8 : data <= 8'hFE;
      10'h1B9 : data <= 8'hC6;
      10'h1BA : data <= 8'h0C;
      10'h1BB : data <= 8'h18;
      10'h1BC : data <= 8'h30;
      10'h1BD : data <= 8'h30;
      10'h1BE : data <= 8'h30;
      10'h1C0 : data <= 8'h7C;
      10'h1C1 : data <= 8'hC6;
      10'h1C2 : data <= 8'hC6;
      10'h1C3 : data <= 8'h7C;
      10'h1C4 : data <= 8'hC6;
      10'h1C5 : data <= 8'hC6;
      10'h1C6 : data <= 8'h7C;
      10'h1C8 : data <= 8'h7C;
      10'h1C9 : data <= 8'hC6;
      10'h1CA : data <= 8'hC6;
      10'h1CB : data <= 8'h7E;
      10'h1CC : data <= 8'h06;
      10'h1CD : data <= 8'h0C;
      10'h1CE : data <= 8'h78;
      10'h1D1 : data <= 8'h18;
      10'h1D2 : data <= 8'h18;
      10'h1D5 : data <= 8'h18;
      10'h1D6 : data <= 8'h18;
      10'h1D9 : data <= 8'h18;
      10'h1DA : data <= 8'h18;
      10'h1DD : data <= 8'h18;
      10'h1DE : data <= 8'h18;
      10'h1DF : data <= 8'h30;
      10'h1E0 : data <= 8'h0C;
      10'h1E1 : data <= 8'h18;
      10'h1E2 : data <= 8'h30;
      10'h1E3 : data <= 8'h60;
      10'h1E4 : data <= 8'h30;
      10'h1E5 : data <= 8'h18;
      10'h1E6 : data <= 8'h0C;
      10'h1EA : data <= 8'h7E;
      10'h1ED : data <= 8'h7E;
      10'h1F0 : data <= 8'h30;
      10'h1F1 : data <= 8'h18;
      10'h1F2 : data <= 8'h0C;
      10'h1F3 : data <= 8'h06;
      10'h1F4 : data <= 8'h0C;
      10'h1F5 : data <= 8'h18;
      10'h1F6 : data <= 8'h30;
      10'h1F8 : data <= 8'h3C;
      10'h1F9 : data <= 8'h66;
      10'h1FA : data <= 8'h06;
      10'h1FB : data <= 8'h0C;
      10'h1FC : data <= 8'h18;
      10'h1FE : data <= 8'h18;
      10'h200 : data <= 8'h7C;
      10'h201 : data <= 8'hC6;
      10'h202 : data <= 8'hDE;
      10'h203 : data <= 8'hDE;
      10'h204 : data <= 8'hDE;
      10'h205 : data <= 8'hC0;
      10'h206 : data <= 8'h7C;
      10'h208 : data <= 8'h38;
      10'h209 : data <= 8'h6C;
      10'h20A : data <= 8'hC6;
      10'h20B : data <= 8'hC6;
      10'h20C : data <= 8'hFE;
      10'h20D : data <= 8'hC6;
      10'h20E : data <= 8'hC6;
      10'h210 : data <= 8'hFC;
      10'h211 : data <= 8'h6E;
      10'h212 : data <= 8'h66;
      10'h213 : data <= 8'h7C;
      10'h214 : data <= 8'h66;
      10'h215 : data <= 8'h6E;
      10'h216 : data <= 8'hFC;
      10'h218 : data <= 8'h3E;
      10'h219 : data <= 8'h62;
      10'h21A : data <= 8'hC0;
      10'h21B : data <= 8'hC0;
      10'h21C : data <= 8'hC0;
      10'h21D : data <= 8'h62;
      10'h21E : data <= 8'h3E;
      10'h220 : data <= 8'hF8;
      10'h221 : data <= 8'h6E;
      10'h222 : data <= 8'h66;
      10'h223 : data <= 8'h66;
      10'h224 : data <= 8'h66;
      10'h225 : data <= 8'h6E;
      10'h226 : data <= 8'hF8;
      10'h228 : data <= 8'hFE;
      10'h229 : data <= 8'h62;
      10'h22A : data <= 8'h60;
      10'h22B : data <= 8'h78;
      10'h22C : data <= 8'h60;
      10'h22D : data <= 8'h62;
      10'h22E : data <= 8'hFE;
      10'h230 : data <= 8'hFE;
      10'h231 : data <= 8'h62;
      10'h232 : data <= 8'h60;
      10'h233 : data <= 8'h78;
      10'h234 : data <= 8'h60;
      10'h235 : data <= 8'h60;
      10'h236 : data <= 8'hF0;
      10'h238 : data <= 8'h3E;
      10'h239 : data <= 8'h62;
      10'h23A : data <= 8'hC0;
      10'h23B : data <= 8'hC0;
      10'h23C : data <= 8'hCE;
      10'h23D : data <= 8'h66;
      10'h23E : data <= 8'h3E;
      10'h240 : data <= 8'hC6;
      10'h241 : data <= 8'hC6;
      10'h242 : data <= 8'hC6;
      10'h243 : data <= 8'hFE;
      10'h244 : data <= 8'hC6;
      10'h245 : data <= 8'hC6;
      10'h246 : data <= 8'hC6;
      10'h248 : data <= 8'h3C;
      10'h249 : data <= 8'h18;
      10'h24A : data <= 8'h18;
      10'h24B : data <= 8'h18;
      10'h24C : data <= 8'h18;
      10'h24D : data <= 8'h18;
      10'h24E : data <= 8'h3C;
      10'h250 : data <= 8'h1E;
      10'h251 : data <= 8'h0C;
      10'h252 : data <= 8'h0C;
      10'h253 : data <= 8'h0C;
      10'h254 : data <= 8'h0C;
      10'h255 : data <= 8'hCC;
      10'h256 : data <= 8'h78;
      10'h258 : data <= 8'hE6;
      10'h259 : data <= 8'h66;
      10'h25A : data <= 8'h6C;
      10'h25B : data <= 8'h78;
      10'h25C : data <= 8'h78;
      10'h25D : data <= 8'h6C;
      10'h25E : data <= 8'hE6;
      10'h260 : data <= 8'hF0;
      10'h261 : data <= 8'h60;
      10'h262 : data <= 8'h60;
      10'h263 : data <= 8'h60;
      10'h264 : data <= 8'h60;
      10'h265 : data <= 8'h66;
      10'h266 : data <= 8'hFE;
      10'h268 : data <= 8'hC6;
      10'h269 : data <= 8'hEE;
      10'h26A : data <= 8'hFE;
      10'h26B : data <= 8'hD6;
      10'h26C : data <= 8'hC6;
      10'h26D : data <= 8'hC6;
      10'h26E : data <= 8'hC6;
      10'h270 : data <= 8'hC6;
      10'h271 : data <= 8'hE6;
      10'h272 : data <= 8'hF6;
      10'h273 : data <= 8'hFE;
      10'h274 : data <= 8'hDE;
      10'h275 : data <= 8'hCE;
      10'h276 : data <= 8'hC6;
      10'h278 : data <= 8'h7C;
      10'h279 : data <= 8'hC6;
      10'h27A : data <= 8'hC6;
      10'h27B : data <= 8'hC6;
      10'h27C : data <= 8'hC6;
      10'h27D : data <= 8'hC6;
      10'h27E : data <= 8'h7C;
      10'h280 : data <= 8'hFC;
      10'h281 : data <= 8'h66;
      10'h282 : data <= 8'h66;
      10'h283 : data <= 8'h7C;
      10'h284 : data <= 8'h60;
      10'h285 : data <= 8'h60;
      10'h286 : data <= 8'hE0;
      10'h288 : data <= 8'h7C;
      10'h289 : data <= 8'hC6;
      10'h28A : data <= 8'hC6;
      10'h28B : data <= 8'hD6;
      10'h28C : data <= 8'hDE;
      10'h28D : data <= 8'h7C;
      10'h28E : data <= 8'h06;
      10'h290 : data <= 8'hFC;
      10'h291 : data <= 8'h66;
      10'h292 : data <= 8'h66;
      10'h293 : data <= 8'h7C;
      10'h294 : data <= 8'h78;
      10'h295 : data <= 8'h6C;
      10'h296 : data <= 8'hE6;
      10'h298 : data <= 8'h7C;
      10'h299 : data <= 8'hC6;
      10'h29A : data <= 8'hE0;
      10'h29B : data <= 8'h38;
      10'h29C : data <= 8'h0E;
      10'h29D : data <= 8'hC6;
      10'h29E : data <= 8'h7C;
      10'h2A0 : data <= 8'h7E;
      10'h2A1 : data <= 8'h5A;
      10'h2A2 : data <= 8'h18;
      10'h2A3 : data <= 8'h18;
      10'h2A4 : data <= 8'h18;
      10'h2A5 : data <= 8'h18;
      10'h2A6 : data <= 8'h3C;
      10'h2A8 : data <= 8'h66;
      10'h2A9 : data <= 8'h66;
      10'h2AA : data <= 8'h66;
      10'h2AB : data <= 8'h66;
      10'h2AC : data <= 8'h66;
      10'h2AD : data <= 8'h66;
      10'h2AE : data <= 8'h3C;
      10'h2B0 : data <= 8'h66;
      10'h2B1 : data <= 8'h66;
      10'h2B2 : data <= 8'h66;
      10'h2B3 : data <= 8'h66;
      10'h2B4 : data <= 8'h66;
      10'h2B5 : data <= 8'h3C;
      10'h2B6 : data <= 8'h18;
      10'h2B8 : data <= 8'hC6;
      10'h2B9 : data <= 8'hC6;
      10'h2BA : data <= 8'hC6;
      10'h2BB : data <= 8'hD6;
      10'h2BC : data <= 8'hFE;
      10'h2BD : data <= 8'hFE;
      10'h2BE : data <= 8'hC6;
      10'h2C0 : data <= 8'hC6;
      10'h2C1 : data <= 8'h6C;
      10'h2C2 : data <= 8'h38;
      10'h2C3 : data <= 8'h38;
      10'h2C4 : data <= 8'h6C;
      10'h2C5 : data <= 8'hC6;
      10'h2C6 : data <= 8'hC6;
      10'h2C8 : data <= 8'h66;
      10'h2C9 : data <= 8'h66;
      10'h2CA : data <= 8'h66;
      10'h2CB : data <= 8'h3C;
      10'h2CC : data <= 8'h18;
      10'h2CD : data <= 8'h18;
      10'h2CE : data <= 8'h3C;
      10'h2D0 : data <= 8'hFE;
      10'h2D1 : data <= 8'hCC;
      10'h2D2 : data <= 8'h18;
      10'h2D3 : data <= 8'h30;
      10'h2D4 : data <= 8'h60;
      10'h2D5 : data <= 8'hC6;
      10'h2D6 : data <= 8'hFE;
      10'h2D8 : data <= 8'h3C;
      10'h2D9 : data <= 8'h30;
      10'h2DA : data <= 8'h30;
      10'h2DB : data <= 8'h30;
      10'h2DC : data <= 8'h30;
      10'h2DD : data <= 8'h30;
      10'h2DE : data <= 8'h3C;
      10'h2E0 : data <= 8'h80;
      10'h2E1 : data <= 8'hC0;
      10'h2E2 : data <= 8'h60;
      10'h2E3 : data <= 8'h30;
      10'h2E4 : data <= 8'h18;
      10'h2E5 : data <= 8'h0C;
      10'h2E6 : data <= 8'h06;
      10'h2E8 : data <= 8'h3C;
      10'h2E9 : data <= 8'h0C;
      10'h2EA : data <= 8'h0C;
      10'h2EB : data <= 8'h0C;
      10'h2EC : data <= 8'h0C;
      10'h2ED : data <= 8'h0C;
      10'h2EE : data <= 8'h3C;
      10'h2F0 : data <= 8'h18;
      10'h2F1 : data <= 8'h3C;
      10'h2F2 : data <= 8'h66;
      10'h2FF : data <= 8'hFF;
      10'h300 : data <= 8'h18;
      10'h301 : data <= 8'h18;
      10'h302 : data <= 8'h0C;
      10'h30A : data <= 8'h38;
      10'h30B : data <= 8'h0C;
      10'h30C : data <= 8'h7C;
      10'h30D : data <= 8'hCC;
      10'h30E : data <= 8'h76;
      10'h310 : data <= 8'h60;
      10'h311 : data <= 8'h60;
      10'h312 : data <= 8'h60;
      10'h313 : data <= 8'h7C;
      10'h314 : data <= 8'h66;
      10'h315 : data <= 8'h66;
      10'h316 : data <= 8'hDC;
      10'h31A : data <= 8'h7C;
      10'h31B : data <= 8'hC4;
      10'h31C : data <= 8'hC0;
      10'h31D : data <= 8'hC4;
      10'h31E : data <= 8'h7C;
      10'h320 : data <= 8'h0C;
      10'h321 : data <= 8'h0C;
      10'h322 : data <= 8'h0C;
      10'h323 : data <= 8'h7C;
      10'h324 : data <= 8'hCC;
      10'h325 : data <= 8'hCC;
      10'h326 : data <= 8'h76;
      10'h32A : data <= 8'h78;
      10'h32B : data <= 8'hCC;
      10'h32C : data <= 8'hFC;
      10'h32D : data <= 8'hC0;
      10'h32E : data <= 8'h7C;
      10'h330 : data <= 8'h38;
      10'h331 : data <= 8'h6C;
      10'h332 : data <= 8'h60;
      10'h333 : data <= 8'hF8;
      10'h334 : data <= 8'h60;
      10'h335 : data <= 8'h60;
      10'h336 : data <= 8'hE0;
      10'h33A : data <= 8'h76;
      10'h33B : data <= 8'hCC;
      10'h33C : data <= 8'hCC;
      10'h33D : data <= 8'h7C;
      10'h33E : data <= 8'h0C;
      10'h33F : data <= 8'h7C;
      10'h340 : data <= 8'hE0;
      10'h341 : data <= 8'h60;
      10'h342 : data <= 8'h60;
      10'h343 : data <= 8'h7C;
      10'h344 : data <= 8'h66;
      10'h345 : data <= 8'h66;
      10'h346 : data <= 8'h66;
      10'h348 : data <= 8'h30;
      10'h34A : data <= 8'h70;
      10'h34B : data <= 8'h30;
      10'h34C : data <= 8'h30;
      10'h34D : data <= 8'h30;
      10'h34E : data <= 8'h38;
      10'h350 : data <= 8'h0C;
      10'h352 : data <= 8'h1C;
      10'h353 : data <= 8'h0C;
      10'h354 : data <= 8'h0C;
      10'h355 : data <= 8'hCC;
      10'h356 : data <= 8'hCC;
      10'h357 : data <= 8'h78;
      10'h358 : data <= 8'hE0;
      10'h359 : data <= 8'h60;
      10'h35A : data <= 8'h66;
      10'h35B : data <= 8'h6C;
      10'h35C : data <= 8'h78;
      10'h35D : data <= 8'h6C;
      10'h35E : data <= 8'h66;
      10'h360 : data <= 8'h70;
      10'h361 : data <= 8'h30;
      10'h362 : data <= 8'h30;
      10'h363 : data <= 8'h30;
      10'h364 : data <= 8'h30;
      10'h365 : data <= 8'h30;
      10'h366 : data <= 8'h38;
      10'h36A : data <= 8'hCC;
      10'h36B : data <= 8'hFE;
      10'h36C : data <= 8'hD6;
      10'h36D : data <= 8'hC6;
      10'h36E : data <= 8'hC6;
      10'h372 : data <= 8'hDC;
      10'h373 : data <= 8'h66;
      10'h374 : data <= 8'h66;
      10'h375 : data <= 8'h66;
      10'h376 : data <= 8'h66;
      10'h37A : data <= 8'h3C;
      10'h37B : data <= 8'h66;
      10'h37C : data <= 8'h66;
      10'h37D : data <= 8'h66;
      10'h37E : data <= 8'h3C;
      10'h382 : data <= 8'hDC;
      10'h383 : data <= 8'h66;
      10'h384 : data <= 8'h66;
      10'h385 : data <= 8'h7C;
      10'h386 : data <= 8'h60;
      10'h387 : data <= 8'hE0;
      10'h38A : data <= 8'h76;
      10'h38B : data <= 8'hCC;
      10'h38C : data <= 8'hCC;
      10'h38D : data <= 8'h7C;
      10'h38E : data <= 8'h0C;
      10'h38F : data <= 8'h0E;
      10'h392 : data <= 8'hDC;
      10'h393 : data <= 8'h76;
      10'h394 : data <= 8'h60;
      10'h395 : data <= 8'h60;
      10'h396 : data <= 8'h60;
      10'h39A : data <= 8'h78;
      10'h39B : data <= 8'hC0;
      10'h39C : data <= 8'h78;
      10'h39D : data <= 8'h0C;
      10'h39E : data <= 8'h78;
      10'h3A0 : data <= 8'h10;
      10'h3A1 : data <= 8'h30;
      10'h3A2 : data <= 8'h78;
      10'h3A3 : data <= 8'h30;
      10'h3A4 : data <= 8'h30;
      10'h3A5 : data <= 8'h34;
      10'h3A6 : data <= 8'h18;
      10'h3AA : data <= 8'hCC;
      10'h3AB : data <= 8'hCC;
      10'h3AC : data <= 8'hCC;
      10'h3AD : data <= 8'hCC;
      10'h3AE : data <= 8'h76;
      10'h3B2 : data <= 8'h66;
      10'h3B3 : data <= 8'h66;
      10'h3B4 : data <= 8'h66;
      10'h3B5 : data <= 8'h3C;
      10'h3B6 : data <= 8'h18;
      10'h3BA : data <= 8'hC6;
      10'h3BB : data <= 8'hC6;
      10'h3BC : data <= 8'hD6;
      10'h3BD : data <= 8'hFE;
      10'h3BE : data <= 8'h6C;
      10'h3C2 : data <= 8'hCC;
      10'h3C3 : data <= 8'h78;
      10'h3C4 : data <= 8'h30;
      10'h3C5 : data <= 8'h78;
      10'h3C6 : data <= 8'hCC;
      10'h3CA : data <= 8'hCC;
      10'h3CB : data <= 8'hCC;
      10'h3CC : data <= 8'hCC;
      10'h3CD : data <= 8'h7C;
      10'h3CE : data <= 8'h0C;
      10'h3CF : data <= 8'h7C;
      10'h3D2 : data <= 8'hFC;
      10'h3D3 : data <= 8'h18;
      10'h3D4 : data <= 8'h30;
      10'h3D5 : data <= 8'h60;
      10'h3D6 : data <= 8'hFC;
      10'h3D8 : data <= 8'h0E;
      10'h3D9 : data <= 8'h18;
      10'h3DA : data <= 8'h18;
      10'h3DB : data <= 8'h70;
      10'h3DC : data <= 8'h18;
      10'h3DD : data <= 8'h18;
      10'h3DE : data <= 8'h0E;
      10'h3E0 : data <= 8'h30;
      10'h3E1 : data <= 8'h30;
      10'h3E2 : data <= 8'h30;
      10'h3E4 : data <= 8'h30;
      10'h3E5 : data <= 8'h30;
      10'h3E6 : data <= 8'h30;
      10'h3E8 : data <= 8'h70;
      10'h3E9 : data <= 8'h18;
      10'h3EA : data <= 8'h18;
      10'h3EB : data <= 8'h0E;
      10'h3EC : data <= 8'h18;
      10'h3ED : data <= 8'h18;
      10'h3EE : data <= 8'h70;
      10'h3F1 : data <= 8'h76;
      10'h3F2 : data <= 8'hDC;
      10'h3F8 : data <= 8'h10;
      10'h3F9 : data <= 8'h38;
      10'h3FA : data <= 8'h6C;
      10'h3FB : data <= 8'hC6;
      10'h3FC : data <= 8'hC6;
      10'h3FD : data <= 8'hC6;
      10'h3FE : data <= 8'hFE;
      default : data <= 8'h00;
    endcase
  end
endmodule
